

	reg signed [9:0] w_r [0:7] = '{9'd256,9'd237,9'd181,9'd98,9'd0,-9'd98,-9'd181,-9'd237};
	reg signed [9:0] w_i [0:7] = '{9'd0,-9'd98,-9'd181,-9'd237,-9'd256,-9'd237,-9'd181,-9'd98};