

	reg signed [9:0] w_r [0:15] = '{9'd256,9'd251,9'd237,9'd213,9'd181,9'd142,9'd98,9'd50,9'd0,-9'd50,-9'd98,-9'd142,-9'd181,-9'd213,-9'd237,-9'd251};
	reg signed [9:0] w_i [0:15] = '{9'd0,-9'd50,-9'd98,-9'd142,-9'd181,-9'd213,-9'd237,-9'd251,-9'd256,-9'd251,-9'd237,-9'd213,-9'd181,-9'd142,-9'd98,-9'd50};