

	reg signed [9:0] w_r [0:3] = '{9'd256,9'd181,9'd0,-9'd181};
	reg signed [9:0] w_i [0:3] = '{9'd0,-9'd181,-9'd256,-9'd181};