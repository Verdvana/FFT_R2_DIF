//=============================================================================
// Module Name:             Butterfly
// Function Description:    FFT butterfly transformation
// Department:              Qualcomm (Shanghai) Co., Ltd.
// Author:                  Verdvana
// Email:                   verdvana@outlook.com
//-----------------------------------------------------------------------------
// Version 	Design		Coding		Simulate    Review      Rel date
// V1.0		Verdvana	Verdvana	Verdvana				2019-11-19
// V2.0		Verdvana	Verdvana	Verdvana				2021-11-21
// V2.1		Verdvana	Verdvana	Verdvana				2021-12-03
//-----------------------------------------------------------------------------
// Version	Modified History
// V1.0		FFT butterfly transformation;
//			DIF;
//			Radix 2;
//			Data width is configurable;
//			The number of sampling points is configurable, BUT the twiddle factor 
//			needs to be calculated in advance and stored in the head file;
//			Pure combinatorial logic.
// V2.0 	Use one stage pipeline design to improve timing;
//			Generate the twiddle factor using the system function, but DC and 
//			Quartus dont support synthesis.
// V2.1		Use a script to generate GENERIC twiddle factors;
//			Twiddle factors are magnified, the magnification needs to be 
//			modified in the script.
//=============================================================================

// Include

// Define
//`define			FPGA_EMU

//Module
module Butterfly #(
	parameter		DATA_WIDTH	= 16,													// Data width
					SERIES 		= 1,													// FFT series
					POW 		= 3     												// The sampling points is N，POW=log2(N)
)(		
	input	wire							clk,										// Clock
	input	wire							rst_n,										// Async reset
	input  	wire	signed [DATA_WIDTH+SERIES*2-1:0]	sink_r [(2)**(POW-SERIES)],		// The real part of the input data
	input  	wire	signed [DATA_WIDTH+SERIES*2-1:0]	sink_i [(2)**(POW-SERIES)],		// The imaginary part of input data
	output 	logic	signed [DATA_WIDTH+SERIES*2+1:0] 	source_r [(2)**(POW-SERIES)],	// The real part of the output data
	output 	logic	signed [DATA_WIDTH+SERIES*2+1:0] 	source_i [(2)**(POW-SERIES)]	// The imaginary part of output data
);

	//=========================================================
	//The time unit and precision of the internal declaration
	timeunit        	1ns;
	timeprecision   	1ps;

    //=========================================================
    // Constant and parameter of twiddle factor
	localparam	GAIN 		= 256,					// Gain of twiddle factor
				N_MAX 		= GAIN*8;				// Maximum sampling points
	localparam int Twiddle_Factor_r [1024] = '{256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,254,254,254,254,254,254,254,254,254,254,253,253,253,253,253,253,253,253,252,252,252,252,252,252,252,252,251,251,251,251,251,251,250,250,250,250,250,250,249,249,249,249,249,249,248,248,248,248,248,247,247,247,247,247,246,246,246,246,245,245,245,245,245,244,244,244,244,243,243,243,243,242,242,242,242,241,241,241,241,240,240,240,239,239,239,239,238,238,238,237,237,237,237,236,236,236,235,235,235,234,234,234,233,233,233,232,232,232,231,231,231,230,230,230,229,229,229,228,228,228,227,227,227,226,226,225,225,225,224,224,224,223,223,222,222,222,221,221,220,220,220,219,219,218,218,218,217,217,216,216,215,215,215,214,214,213,213,212,212,212,211,211,210,210,209,209,208,208,207,207,207,206,206,205,205,204,204,203,203,202,202,201,201,200,200,199,199,198,198,197,197,196,196,195,195,194,194,193,193,192,192,191,191,190,190,189,189,188,188,187,186,186,185,185,184,184,183,183,182,182,181,180,180,179,179,178,178,177,177,176,175,175,174,174,173,173,172,171,171,170,170,169,168,168,167,167,166,165,165,164,164,163,162,162,161,161,160,159,159,158,158,157,156,156,155,154,154,153,153,152,151,151,150,149,149,148,147,147,146,145,145,144,144,143,142,142,141,140,140,139,138,138,137,136,136,135,134,134,133,132,132,131,130,130,129,128,128,127,126,126,125,124,123,123,122,121,121,120,119,119,118,117,117,116,115,114,114,113,112,112,111,110,109,109,108,107,107,106,105,104,104,103,102,102,101,100,99,99,98,97,97,96,95,94,94,93,92,91,91,90,89,88,88,87,86,86,85,84,83,83,82,81,80,80,79,78,77,77,76,75,74,74,73,72,71,71,70,69,68,68,67,66,65,64,64,63,62,61,61,60,59,58,58,57,56,55,55,54,53,52,51,51,50,49,48,48,47,46,45,45,44,43,42,41,41,40,39,38,38,37,36,35,34,34,33,32,31,31,30,29,28,27,27,26,25,24,24,23,22,21,20,20,19,18,17,16,16,15,14,13,13,12,11,10,9,9,8,7,6,6,5,4,3,2,2,1,0,-1,-2,-2,-3,-4,-5,-5,-6,-7,-8,-9,-9,-10,-11,-12,-13,-13,-14,-15,-16,-16,-17,-18,-19,-20,-20,-21,-22,-23,-24,-24,-25,-26,-27,-27,-28,-29,-30,-31,-31,-32,-33,-34,-34,-35,-36,-37,-38,-38,-39,-40,-41,-41,-42,-43,-44,-45,-45,-46,-47,-48,-48,-49,-50,-51,-51,-52,-53,-54,-55,-55,-56,-57,-58,-58,-59,-60,-61,-61,-62,-63,-64,-64,-65,-66,-67,-68,-68,-69,-70,-71,-71,-72,-73,-74,-74,-75,-76,-77,-77,-78,-79,-80,-80,-81,-82,-83,-83,-84,-85,-85,-86,-87,-88,-88,-89,-90,-91,-91,-92,-93,-94,-94,-95,-96,-97,-97,-98,-99,-99,-100,-101,-102,-102,-103,-104,-104,-105,-106,-107,-107,-108,-109,-109,-110,-111,-112,-112,-113,-114,-114,-115,-116,-116,-117,-118,-119,-119,-120,-121,-121,-122,-123,-123,-124,-125,-125,-126,-127,-128,-128,-129,-130,-130,-131,-132,-132,-133,-134,-134,-135,-136,-136,-137,-138,-138,-139,-140,-140,-141,-142,-142,-143,-144,-144,-145,-145,-146,-147,-147,-148,-149,-149,-150,-151,-151,-152,-152,-153,-154,-154,-155,-156,-156,-157,-157,-158,-159,-159,-160,-161,-161,-162,-162,-163,-164,-164,-165,-165,-166,-167,-167,-168,-168,-169,-170,-170,-171,-171,-172,-172,-173,-174,-174,-175,-175,-176,-177,-177,-178,-178,-179,-179,-180,-180,-181,-182,-182,-183,-183,-184,-184,-185,-185,-186,-186,-187,-188,-188,-189,-189,-190,-190,-191,-191,-192,-192,-193,-193,-194,-194,-195,-195,-196,-196,-197,-197,-198,-198,-199,-199,-200,-200,-201,-201,-202,-202,-203,-203,-204,-204,-205,-205,-206,-206,-207,-207,-207,-208,-208,-209,-209,-210,-210,-211,-211,-212,-212,-212,-213,-213,-214,-214,-215,-215,-215,-216,-216,-217,-217,-218,-218,-218,-219,-219,-220,-220,-220,-221,-221,-222,-222,-222,-223,-223,-224,-224,-224,-225,-225,-225,-226,-226,-226,-227,-227,-228,-228,-228,-229,-229,-229,-230,-230,-230,-231,-231,-231,-232,-232,-232,-233,-233,-233,-234,-234,-234,-235,-235,-235,-236,-236,-236,-237,-237,-237,-237,-238,-238,-238,-239,-239,-239,-239,-240,-240,-240,-240,-241,-241,-241,-242,-242,-242,-242,-243,-243,-243,-243,-244,-244,-244,-244,-245,-245,-245,-245,-245,-246,-246,-246,-246,-247,-247,-247,-247,-247,-248,-248,-248,-248,-248,-249,-249,-249,-249,-249,-249,-250,-250,-250,-250,-250,-250,-251,-251,-251,-251,-251,-251,-252,-252,-252,-252,-252,-252,-252,-252,-253,-253,-253,-253,-253,-253,-253,-253,-254,-254,-254,-254,-254,-254,-254,-254,-254,-254,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256};
	localparam int Twiddle_Factor_i [1024] = '{0,-1,-2,-2,-3,-4,-5,-5,-6,-7,-8,-9,-9,-10,-11,-12,-13,-13,-14,-15,-16,-16,-17,-18,-19,-20,-20,-21,-22,-23,-24,-24,-25,-26,-27,-27,-28,-29,-30,-31,-31,-32,-33,-34,-34,-35,-36,-37,-38,-38,-39,-40,-41,-41,-42,-43,-44,-45,-45,-46,-47,-48,-48,-49,-50,-51,-51,-52,-53,-54,-55,-55,-56,-57,-58,-58,-59,-60,-61,-61,-62,-63,-64,-64,-65,-66,-67,-68,-68,-69,-70,-71,-71,-72,-73,-74,-74,-75,-76,-77,-77,-78,-79,-80,-80,-81,-82,-83,-83,-84,-85,-86,-86,-87,-88,-88,-89,-90,-91,-91,-92,-93,-94,-94,-95,-96,-97,-97,-98,-99,-99,-100,-101,-102,-102,-103,-104,-104,-105,-106,-107,-107,-108,-109,-109,-110,-111,-112,-112,-113,-114,-114,-115,-116,-116,-117,-118,-119,-119,-120,-121,-121,-122,-123,-123,-124,-125,-125,-126,-127,-128,-128,-129,-130,-130,-131,-132,-132,-133,-134,-134,-135,-136,-136,-137,-138,-138,-139,-140,-140,-141,-142,-142,-143,-144,-144,-145,-145,-146,-147,-147,-148,-149,-149,-150,-151,-151,-152,-152,-153,-154,-154,-155,-156,-156,-157,-157,-158,-159,-159,-160,-161,-161,-162,-162,-163,-164,-164,-165,-165,-166,-167,-167,-168,-168,-169,-170,-170,-171,-171,-172,-172,-173,-174,-174,-175,-175,-176,-177,-177,-178,-178,-179,-179,-180,-180,-181,-182,-182,-183,-183,-184,-184,-185,-185,-186,-186,-187,-188,-188,-189,-189,-190,-190,-191,-191,-192,-192,-193,-193,-194,-194,-195,-195,-196,-196,-197,-197,-198,-198,-199,-199,-200,-200,-201,-201,-202,-202,-203,-203,-204,-204,-205,-205,-206,-206,-207,-207,-207,-208,-208,-209,-209,-210,-210,-211,-211,-212,-212,-212,-213,-213,-214,-214,-215,-215,-215,-216,-216,-217,-217,-218,-218,-218,-219,-219,-220,-220,-220,-221,-221,-222,-222,-222,-223,-223,-224,-224,-224,-225,-225,-225,-226,-226,-227,-227,-227,-228,-228,-228,-229,-229,-229,-230,-230,-230,-231,-231,-231,-232,-232,-232,-233,-233,-233,-234,-234,-234,-235,-235,-235,-236,-236,-236,-237,-237,-237,-237,-238,-238,-238,-239,-239,-239,-239,-240,-240,-240,-240,-241,-241,-241,-242,-242,-242,-242,-243,-243,-243,-243,-244,-244,-244,-244,-245,-245,-245,-245,-245,-246,-246,-246,-246,-247,-247,-247,-247,-247,-248,-248,-248,-248,-248,-249,-249,-249,-249,-249,-249,-250,-250,-250,-250,-250,-250,-251,-251,-251,-251,-251,-251,-252,-252,-252,-252,-252,-252,-252,-252,-253,-253,-253,-253,-253,-253,-253,-253,-254,-254,-254,-254,-254,-254,-254,-254,-254,-254,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-256,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-255,-254,-254,-254,-254,-254,-254,-254,-254,-254,-254,-253,-253,-253,-253,-253,-253,-253,-253,-252,-252,-252,-252,-252,-252,-252,-252,-251,-251,-251,-251,-251,-251,-250,-250,-250,-250,-250,-250,-249,-249,-249,-249,-249,-249,-248,-248,-248,-248,-248,-247,-247,-247,-247,-247,-246,-246,-246,-246,-245,-245,-245,-245,-245,-244,-244,-244,-244,-243,-243,-243,-243,-242,-242,-242,-242,-241,-241,-241,-241,-240,-240,-240,-239,-239,-239,-239,-238,-238,-238,-237,-237,-237,-237,-236,-236,-236,-235,-235,-235,-234,-234,-234,-233,-233,-233,-232,-232,-232,-231,-231,-231,-230,-230,-230,-229,-229,-229,-228,-228,-228,-227,-227,-227,-226,-226,-225,-225,-225,-224,-224,-224,-223,-223,-222,-222,-222,-221,-221,-220,-220,-220,-219,-219,-218,-218,-218,-217,-217,-216,-216,-215,-215,-215,-214,-214,-213,-213,-212,-212,-212,-211,-211,-210,-210,-209,-209,-208,-208,-207,-207,-207,-206,-206,-205,-205,-204,-204,-203,-203,-202,-202,-201,-201,-200,-200,-199,-199,-198,-198,-197,-197,-196,-196,-195,-195,-194,-194,-193,-193,-192,-192,-191,-191,-190,-190,-189,-189,-188,-188,-187,-186,-186,-185,-185,-184,-184,-183,-183,-182,-182,-181,-180,-180,-179,-179,-178,-178,-177,-177,-176,-175,-175,-174,-174,-173,-173,-172,-171,-171,-170,-170,-169,-168,-168,-167,-167,-166,-165,-165,-164,-164,-163,-162,-162,-161,-161,-160,-159,-159,-158,-158,-157,-156,-156,-155,-154,-154,-153,-153,-152,-151,-151,-150,-149,-149,-148,-147,-147,-146,-145,-145,-144,-144,-143,-142,-142,-141,-140,-140,-139,-138,-138,-137,-136,-136,-135,-134,-134,-133,-132,-132,-131,-130,-130,-129,-128,-128,-127,-126,-126,-125,-124,-123,-123,-122,-121,-121,-120,-119,-119,-118,-117,-117,-116,-115,-114,-114,-113,-112,-112,-111,-110,-109,-109,-108,-107,-107,-106,-105,-104,-104,-103,-102,-102,-101,-100,-99,-99,-98,-97,-97,-96,-95,-94,-94,-93,-92,-91,-91,-90,-89,-88,-88,-87,-86,-86,-85,-84,-83,-83,-82,-81,-80,-80,-79,-78,-77,-77,-76,-75,-74,-74,-73,-72,-71,-71,-70,-69,-68,-68,-67,-66,-65,-65,-64,-63,-62,-61,-61,-60,-59,-58,-58,-57,-56,-55,-55,-54,-53,-52,-52,-51,-50,-49,-48,-48,-47,-46,-45,-45,-44,-43,-42,-41,-41,-40,-39,-38,-38,-37,-36,-35,-34,-34,-33,-32,-31,-31,-30,-29,-28,-27,-27,-26,-25,-24,-24,-23,-22,-21,-20,-20,-19,-18,-17,-17,-16,-15,-14,-13,-13,-12,-11,-10,-9,-9,-8,-7,-6,-6,-5,-4,-3,-2,-2,-1};

    //=========================================================
    // Local parameter
    localparam 	DATA_NUM 	= 2**(POW-SERIES),		// Data number
				SHIFT_L		= $clog2(GAIN),			// Bits of left shifts
				TCO			= 0.2;					// Simulate the delay of the register
    //=========================================================
    // Function
    /* DC and Quartus dont support synthesis the following system functions like "$cos $sin", but Vivado do. Is very smart!
	function shortint Twiddle_Factor_r;
	input int i;
		Twiddle_Factor_r = $cos( 2*3.1415*(i/((2**POW)/DATA_NUM)))*GAIN;
	endfunction
	function shortint Twiddle_Factor_i;
	input int i;
		Twiddle_Factor_i = $sin(-2*3.1415*(i/((2**POW)/DATA_NUM)))*GAIN;
	endfunction
    */

    //=========================================================
	// The first half of the butterfly transformation
    logic signed [DATA_WIDTH+SERIES*2+1:0]	sum_re [DATA_NUM/2];
    logic signed [DATA_WIDTH+SERIES*2+1:0]	sum_im [DATA_NUM/2];

    always_ff@(posedge clk, negedge rst_n) begin
        if(!rst_n)
            for(int i=0;i<(DATA_NUM/2);i++)begin
                sum_re[i]	<= #TCO '0;
                sum_im[i]	<= #TCO '0;
            end
        else
            for(int i=0;i<(DATA_NUM/2);i++)begin
                sum_re[i]	<= #TCO ( sink_r[i] + sink_r[i+DATA_NUM/2] );
                sum_im[i]	<= #TCO ( sink_i[i] + sink_i[i+DATA_NUM/2] );
            end
    end

	always_ff@(posedge clk, negedge rst_n)begin
		if(!rst_n)
			for(int i=0;i<(DATA_NUM/2);i++)begin
				source_r[i]	<= #TCO '0;
				source_i[i]	<= #TCO '0;
			end
		else
			for(int i=0;i<(DATA_NUM/2);i++)begin
				source_r[i]	<= #TCO sum_re[i];
				source_i[i]	<= #TCO sum_im[i];
			end
	end


	//====================================================
	// The second half of the butterfly transformation
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2:0]	product_re_1	[DATA_NUM/2];	// Product of real
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2:0]	product_re_2	[DATA_NUM/2];
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2:0]	product_im_1	[DATA_NUM/2];	// Product of imaginary
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2:0]	product_im_2	[DATA_NUM/2];
    
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2+1:0]	plural_re		[DATA_NUM/2];	// Result of real
	logic signed [DATA_WIDTH+SHIFT_L+SERIES*2+1:0]	plural_im		[DATA_NUM/2];	// Result of imaginary

	always_ff@(posedge clk, negedge rst_n)begin
        if(!rst_n)
            for(int i=(DATA_NUM/2);i<DATA_NUM;i++)begin
                product_re_1[i-DATA_NUM/2]	<= #TCO '0;
				product_re_2[i-DATA_NUM/2]	<= #TCO '0;

				product_im_1[i-DATA_NUM/2]	<= #TCO '0;
				product_im_2[i-DATA_NUM/2]	<= #TCO '0;
            end
        else
			for(int i=(DATA_NUM/2);i<DATA_NUM;i++)begin
			    product_re_1[i-DATA_NUM/2]	<= #TCO ( sink_r[i-DATA_NUM/2] - sink_r[i] ) * Twiddle_Factor_r[(i-DATA_NUM/2)*N_MAX/DATA_NUM];	//Before simplify: Twiddle_Factor_r[(i-DATA_NUM/2)*((2**POW)/DATA_NUM) * (N_MAX/(2**POW))]
			    product_re_2[i-DATA_NUM/2]	<= #TCO ( sink_i[i-DATA_NUM/2] - sink_i[i] ) * Twiddle_Factor_i[(i-DATA_NUM/2)*N_MAX/DATA_NUM];

			    product_im_1[i-DATA_NUM/2]	<= #TCO ( sink_r[i-DATA_NUM/2] - sink_r[i] ) * Twiddle_Factor_i[(i-DATA_NUM/2)*N_MAX/DATA_NUM];
			    product_im_2[i-DATA_NUM/2]	<= #TCO ( sink_i[i-DATA_NUM/2] - sink_i[i] ) * Twiddle_Factor_r[(i-DATA_NUM/2)*N_MAX/DATA_NUM];
			end
	end

    always_comb begin
        for(int i=(DATA_NUM/2);i<DATA_NUM;i++)begin
            plural_re[i-DATA_NUM/2]	= product_re_1[i-DATA_NUM/2] - product_re_2[i-DATA_NUM/2];
            plural_im[i-DATA_NUM/2]	= product_im_1[i-DATA_NUM/2] + product_im_2[i-DATA_NUM/2];
        end
    end

	always_ff@(posedge clk, negedge rst_n)begin
		if(!rst_n)
			for(int i=(DATA_NUM/2);i<DATA_NUM;i++)begin
				source_r[i]	<= #TCO '0;
				source_i[i]	<= #TCO '0;
			end
		else
			for(int i=(DATA_NUM/2);i<DATA_NUM;i++)begin
				source_r[i]	<= #TCO plural_re[i-DATA_NUM/2] >>> SHIFT_L;
				source_i[i]	<= #TCO plural_im[i-DATA_NUM/2] >>> SHIFT_L;
			end
	end

endmodule
