	reg signed [9:0] w_r [0:31] = '{9'd256,9'd255,9'd251,9'd245,9'd237,9'd226,9'd213,9'd198,9'd181,9'd162,9'd142,9'd121,9'd98,9'd74,9'd50,9'd25,9'd0,-9'd25,-9'd50,-9'd74,-9'd98,-9'd121,-9'd142,-9'd162,-9'd181,-9'd198,-9'd213,-9'd226,-9'd237,-9'd245,-9'd251,-9'd255};
	reg signed [9:0] w_i [0:31] = '{9'd0,-9'd25,-9'd50,-9'd74,-9'd98,-9'd121,-9'd142,-9'd162,-9'd181,-9'd198,-9'd213,-9'd226,-9'd237,-9'd245,-9'd251,-9'd255,-9'd256,-9'd255,-9'd251,-9'd245,-9'd237,-9'd226,-9'd213,-9'd198,-9'd181,-9'd162,-9'd142,-9'd121,-9'd98,-9'd74,-9'd50,-9'd25};